library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity full_adder is 
	port(bit1 : in std_logic;
	     bit2 : in std_logic;
	     cin  : in std_logic;
	     S : out std_logic;	-- sum
	     C : out std_logic); -- carry
end full_adder;

architecture fullAdderLogic of full_adder is
component half_adder is
port(bit1 : in std_logic;
     bit2 : in std_logic;
     S : out std_logic;	-- sum
     C : out std_logic); -- carry
end component;

signal C1, C2, S1 : std_logic;

begin 
ha1: half_adder
	port map (bit1, bit2, S1, C1);
ha2: half_adder 
	port map (S1, cin, S, C2);
C <= C1 or C2;
end fullAdderLogic;
